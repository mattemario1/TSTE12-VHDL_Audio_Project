--
-- VHDL Architecture The_Reverb_Revolutionary_lib.graphic_gen.graphic_gen_arch
--
-- Created:
--          by - emipi270.student-liu.se (muxen2-114.ad.liu.se)
--          at - 13:34:19 10/02/24
--
-- using Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 18:06:06
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY Visual_graphic_gen IS
-- Declarations

END Visual_graphic_gen ;

--
ARCHITECTURE graphic_gen_arch OF Visual_graphic_gen IS
BEGIN
END ARCHITECTURE graphic_gen_arch;










