
--
ARCHITECTURE Group_no_arch OF Group_no_ent IS
BEGIN
  
  HEX7 <= "1000000"; --0
  HEX6 <= "0010010"; --5
  
END ARCHITECTURE Group_no_arch;

